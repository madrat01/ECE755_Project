package defines_pkg;
    typedef enum logic [1:0] {IDLE, DNN0_DNN1_Y_OUT, DNN2_DNN3_Y_OUT, FINAL_OUT} dnn_state_t;
endpackage
